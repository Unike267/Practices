-- #################################################################################################
-- # << NEORV32 - Test Setup using the default UART-Bootloader to upload and run executables >>    #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # The NEORV32 RISC-V Processor - https://github.com/stnolting/neorv32                           #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library neorv32;
use neorv32.neorv32_package.all;

entity neorv32_multp_wishbone is
  generic (
    -- adapt these for your setup --
    CLOCK_FREQUENCY   : natural := 100000000; -- clock frequency of clk_i in Hz
    MEM_INT_IMEM_SIZE : natural := 6*1024;   -- size of processor-internal instruction memory in bytes
    MEM_INT_DMEM_SIZE : natural := 8*1024     -- size of processor-internal data memory in bytes
  );
  port (
    -- Global control --
    clk_i       : in  std_ulogic; -- global clock, rising edge
    rstn_i      : in  std_ulogic; -- global reset, low-active, async
    -- GPIO --
    gpio_o      : out std_ulogic_vector(7 downto 0); -- parallel output
    -- UART0 --
    uart0_txd_o : out std_ulogic; -- UART0 send data
    uart0_rxd_i : in  std_ulogic  -- UART0 receive data
  );
end entity;

architecture neorv32_multp_wishbone_rtl of neorv32_multp_wishbone is

  signal con_gpio_o : std_ulogic_vector(63 downto 0);

-- Declaration of mult_wrapper axi buffer constants

constant N_bits : natural := 32; -- 32 bits (16 bits plus 16 bits)

-- Declaration of wishbone signals

signal wb_we_o : std_logic;
signal wb_stb_o : std_logic;
signal wb_ack_i : std_logic;
signal wb_cyc_o : std_logic;
signal wb_err_i : std_logic;

signal wb_adr_o : std_logic_vector(31 downto 0);
signal wb_dat_i : std_logic_vector(31 downto 0);
signal wb_dat_o : std_logic_vector(31 downto 0);
signal wb_sel_o : std_logic_vector(3 downto 0);

signal wb_adr_o_u : std_ulogic_vector(31 downto 0);
signal wb_dat_i_u : std_ulogic_vector(31 downto 0);
signal wb_dat_o_u : std_ulogic_vector(31 downto 0);
signal wb_sel_o_u : std_ulogic_vector(3 downto 0);

-- Signals for debug
--attribute MARK_DEBUG : string;
--attribute MARK_DEBUG of wb_stb_o,wb_cyc_o,wb_ack_i,wb_adr_o,wb_dat_i,wb_dat_o,wb_sel_o : signal is "true";

begin

-- Multp wishbone wrapper instantation

multp_wishbone_0 : entity work.multp_wishbone
                                generic map(  
                                        N_bits => N_bits
                                        )
                                port map(
                                    rst_i => rstn_i,
                                    clk_i => clk_i,
                                    adr_i => wb_adr_o,
                                    dat_i => wb_dat_o,
                                    dat_o => wb_dat_i,
                                    we_i => wb_we_o,
                                    sel_i => wb_sel_o,
                                    stb_i => wb_stb_o,
                                    ack_o => wb_ack_i,
                                    cyc_i => wb_cyc_o,
                                    err_o => wb_err_i,
                                    stall_o => open
                                    );

  -- The Core Of The Problem ----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_top_inst: neorv32_top
  generic map (
    -- General --
    CLOCK_FREQUENCY              => CLOCK_FREQUENCY,   -- clock frequency of clk_i in Hz
    INT_BOOTLOADER_EN            => false,              -- boot configuration: true = boot explicit bootloader; false = boot from int/ext (I)MEM
    -- RISC-V CPU Extensions --
    CPU_EXTENSION_RISCV_C        => true,              -- implement compressed extension?
    CPU_EXTENSION_RISCV_M        => true,              -- implement mul/div extension?
    CPU_EXTENSION_RISCV_Zicntr   => true,              -- implement base counters?
    -- Internal Instruction memory --
    MEM_INT_IMEM_EN              => true,              -- implement processor-internal instruction memory
    MEM_INT_IMEM_SIZE            => MEM_INT_IMEM_SIZE, -- size of processor-internal instruction memory in bytes
    -- Internal Data memory --
    MEM_INT_DMEM_EN              => true,              -- implement processor-internal data memory
    MEM_INT_DMEM_SIZE            => MEM_INT_DMEM_SIZE, -- size of processor-internal data memory in bytes
    -- Processor peripherals --
    IO_GPIO_NUM                  => 8,                 -- number of GPIO input/output pairs (0..64)
    IO_MTIME_EN                  => true,              -- implement machine system timer (MTIME)?
    IO_UART0_EN                  => true,              -- implement primary universal asynchronous receiver/transmitter (UART0)?
    -- XBUS (WISHBONE) --
    XBUS_EN                      => true,              -- implement XBUS interface?
    XBUS_TIMEOUT                 => 4096,              -- cycles after a pending bus access auto-terminates (0 = disabled)
    XBUS_REGSTAGE_EN             => false,             -- add XBUS register stage
    XBUS_CACHE_EN                => false              -- enable external bus cache (x-cache)
  )
  port map (
    -- Global control --
    clk_i       => clk_i,       -- global clock, rising edge
    rstn_i      => rstn_i,      -- global reset, low-active, async
    -- GPIO (available if IO_GPIO_EN = true) --
    gpio_o      => con_gpio_o,  -- parallel output
    -- primary UART0 (available if IO_GPIO_NUM > 0) --
    uart0_txd_o => uart0_txd_o, -- UART0 send data
    uart0_rxd_i => uart0_rxd_i,  -- UART0 receive data
    -- Wishbone (XBUS) interface --
    xbus_adr_o    => wb_adr_o_u,    -- address
    xbus_dat_i    => wb_dat_i_u,    -- read data
    xbus_dat_o    => wb_dat_o_u,    -- write data
    xbus_we_o     => wb_we_o,     -- read/write
    xbus_sel_o    => wb_sel_o_u,    -- byte enable
    xbus_stb_o    => wb_stb_o,    -- strobe
    xbus_cyc_o    => wb_cyc_o,    -- valid cycle
    xbus_ack_i    => wb_ack_i,    -- transfer acknowledge
    xbus_err_i    => wb_err_i     -- transfer error
  );

-- GPIO output --
gpio_o <= con_gpio_o(7 downto 0);

-- Adjust with ulogic:

wb_adr_o <= To_StdLogicVector(wb_adr_o_u);
wb_dat_o <= To_StdLogicVector(wb_dat_o_u);
wb_sel_o <= To_StdLogicVector(wb_sel_o_u);

wb_dat_i_u <= To_StdULogicVector(wb_dat_i);

end architecture;

